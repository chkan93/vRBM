`define TEST_BENCH
`include "../config.v"
`include "../RBMLayer.v"


module test_RBMLayer;



endmodule

`define TEST_BENCH
`include "../config.v"
`include "../ClassifyLayer.v"


module test_ClassifyLayer;



endmodule
